##
## LEF for PtnCells ;
## created by Innovus v18.10-p002_1 on Wed Mar 31 16:31:48 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO aes128key
  CLASS BLOCK ;
  SIZE 251.180000 BY 248.920000 ;
  FOREIGN aes128key 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.290000 248.850000 3.360000 248.920000 ;
    END
  END reset
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
  END clock
  PIN empty
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 248.200000 0.000000 248.270000 0.070000 ;
    END
  END empty
  PIN load
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 4.240000 248.850000 4.310000 248.920000 ;
    END
  END load
  PIN key[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 125.840000 248.850000 125.910000 248.920000 ;
    END
  END key[127]
  PIN key[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 124.890000 248.850000 124.960000 248.920000 ;
    END
  END key[126]
  PIN key[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 123.940000 248.850000 124.010000 248.920000 ;
    END
  END key[125]
  PIN key[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 122.990000 248.850000 123.060000 248.920000 ;
    END
  END key[124]
  PIN key[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 122.040000 248.850000 122.110000 248.920000 ;
    END
  END key[123]
  PIN key[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.090000 248.850000 121.160000 248.920000 ;
    END
  END key[122]
  PIN key[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 120.140000 248.850000 120.210000 248.920000 ;
    END
  END key[121]
  PIN key[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 119.190000 248.850000 119.260000 248.920000 ;
    END
  END key[120]
  PIN key[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 118.240000 248.850000 118.310000 248.920000 ;
    END
  END key[119]
  PIN key[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 117.290000 248.850000 117.360000 248.920000 ;
    END
  END key[118]
  PIN key[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 116.340000 248.850000 116.410000 248.920000 ;
    END
  END key[117]
  PIN key[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 115.390000 248.850000 115.460000 248.920000 ;
    END
  END key[116]
  PIN key[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 114.440000 248.850000 114.510000 248.920000 ;
    END
  END key[115]
  PIN key[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 113.490000 248.850000 113.560000 248.920000 ;
    END
  END key[114]
  PIN key[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 112.540000 248.850000 112.610000 248.920000 ;
    END
  END key[113]
  PIN key[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 111.590000 248.850000 111.660000 248.920000 ;
    END
  END key[112]
  PIN key[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 110.640000 248.850000 110.710000 248.920000 ;
    END
  END key[111]
  PIN key[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 109.690000 248.850000 109.760000 248.920000 ;
    END
  END key[110]
  PIN key[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 108.740000 248.850000 108.810000 248.920000 ;
    END
  END key[109]
  PIN key[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 107.790000 248.850000 107.860000 248.920000 ;
    END
  END key[108]
  PIN key[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 106.840000 248.850000 106.910000 248.920000 ;
    END
  END key[107]
  PIN key[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 105.890000 248.850000 105.960000 248.920000 ;
    END
  END key[106]
  PIN key[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 104.940000 248.850000 105.010000 248.920000 ;
    END
  END key[105]
  PIN key[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 103.990000 248.850000 104.060000 248.920000 ;
    END
  END key[104]
  PIN key[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 103.040000 248.850000 103.110000 248.920000 ;
    END
  END key[103]
  PIN key[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 102.090000 248.850000 102.160000 248.920000 ;
    END
  END key[102]
  PIN key[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 101.140000 248.850000 101.210000 248.920000 ;
    END
  END key[101]
  PIN key[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 100.190000 248.850000 100.260000 248.920000 ;
    END
  END key[100]
  PIN key[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 99.240000 248.850000 99.310000 248.920000 ;
    END
  END key[99]
  PIN key[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 98.290000 248.850000 98.360000 248.920000 ;
    END
  END key[98]
  PIN key[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 97.340000 248.850000 97.410000 248.920000 ;
    END
  END key[97]
  PIN key[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 96.390000 248.850000 96.460000 248.920000 ;
    END
  END key[96]
  PIN key[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 95.440000 248.850000 95.510000 248.920000 ;
    END
  END key[95]
  PIN key[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 94.490000 248.850000 94.560000 248.920000 ;
    END
  END key[94]
  PIN key[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 93.540000 248.850000 93.610000 248.920000 ;
    END
  END key[93]
  PIN key[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 92.590000 248.850000 92.660000 248.920000 ;
    END
  END key[92]
  PIN key[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 91.640000 248.850000 91.710000 248.920000 ;
    END
  END key[91]
  PIN key[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 90.690000 248.850000 90.760000 248.920000 ;
    END
  END key[90]
  PIN key[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 89.740000 248.850000 89.810000 248.920000 ;
    END
  END key[89]
  PIN key[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 88.790000 248.850000 88.860000 248.920000 ;
    END
  END key[88]
  PIN key[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 87.840000 248.850000 87.910000 248.920000 ;
    END
  END key[87]
  PIN key[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 86.890000 248.850000 86.960000 248.920000 ;
    END
  END key[86]
  PIN key[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 85.940000 248.850000 86.010000 248.920000 ;
    END
  END key[85]
  PIN key[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 84.990000 248.850000 85.060000 248.920000 ;
    END
  END key[84]
  PIN key[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 84.040000 248.850000 84.110000 248.920000 ;
    END
  END key[83]
  PIN key[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 83.090000 248.850000 83.160000 248.920000 ;
    END
  END key[82]
  PIN key[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 82.140000 248.850000 82.210000 248.920000 ;
    END
  END key[81]
  PIN key[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 81.190000 248.850000 81.260000 248.920000 ;
    END
  END key[80]
  PIN key[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 80.240000 248.850000 80.310000 248.920000 ;
    END
  END key[79]
  PIN key[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 79.290000 248.850000 79.360000 248.920000 ;
    END
  END key[78]
  PIN key[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 78.340000 248.850000 78.410000 248.920000 ;
    END
  END key[77]
  PIN key[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 77.390000 248.850000 77.460000 248.920000 ;
    END
  END key[76]
  PIN key[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 76.440000 248.850000 76.510000 248.920000 ;
    END
  END key[75]
  PIN key[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 75.490000 248.850000 75.560000 248.920000 ;
    END
  END key[74]
  PIN key[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 74.540000 248.850000 74.610000 248.920000 ;
    END
  END key[73]
  PIN key[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 73.590000 248.850000 73.660000 248.920000 ;
    END
  END key[72]
  PIN key[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 72.640000 248.850000 72.710000 248.920000 ;
    END
  END key[71]
  PIN key[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 71.690000 248.850000 71.760000 248.920000 ;
    END
  END key[70]
  PIN key[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 70.740000 248.850000 70.810000 248.920000 ;
    END
  END key[69]
  PIN key[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 69.790000 248.850000 69.860000 248.920000 ;
    END
  END key[68]
  PIN key[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 68.840000 248.850000 68.910000 248.920000 ;
    END
  END key[67]
  PIN key[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 67.890000 248.850000 67.960000 248.920000 ;
    END
  END key[66]
  PIN key[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 66.940000 248.850000 67.010000 248.920000 ;
    END
  END key[65]
  PIN key[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 65.990000 248.850000 66.060000 248.920000 ;
    END
  END key[64]
  PIN key[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 65.040000 248.850000 65.110000 248.920000 ;
    END
  END key[63]
  PIN key[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 64.090000 248.850000 64.160000 248.920000 ;
    END
  END key[62]
  PIN key[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 63.140000 248.850000 63.210000 248.920000 ;
    END
  END key[61]
  PIN key[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 62.190000 248.850000 62.260000 248.920000 ;
    END
  END key[60]
  PIN key[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 61.240000 248.850000 61.310000 248.920000 ;
    END
  END key[59]
  PIN key[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 60.290000 248.850000 60.360000 248.920000 ;
    END
  END key[58]
  PIN key[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 59.340000 248.850000 59.410000 248.920000 ;
    END
  END key[57]
  PIN key[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 58.390000 248.850000 58.460000 248.920000 ;
    END
  END key[56]
  PIN key[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 57.440000 248.850000 57.510000 248.920000 ;
    END
  END key[55]
  PIN key[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 56.490000 248.850000 56.560000 248.920000 ;
    END
  END key[54]
  PIN key[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 55.540000 248.850000 55.610000 248.920000 ;
    END
  END key[53]
  PIN key[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 54.590000 248.850000 54.660000 248.920000 ;
    END
  END key[52]
  PIN key[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 53.640000 248.850000 53.710000 248.920000 ;
    END
  END key[51]
  PIN key[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 52.690000 248.850000 52.760000 248.920000 ;
    END
  END key[50]
  PIN key[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 51.740000 248.850000 51.810000 248.920000 ;
    END
  END key[49]
  PIN key[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 50.790000 248.850000 50.860000 248.920000 ;
    END
  END key[48]
  PIN key[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 49.840000 248.850000 49.910000 248.920000 ;
    END
  END key[47]
  PIN key[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 48.890000 248.850000 48.960000 248.920000 ;
    END
  END key[46]
  PIN key[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 47.940000 248.850000 48.010000 248.920000 ;
    END
  END key[45]
  PIN key[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 46.990000 248.850000 47.060000 248.920000 ;
    END
  END key[44]
  PIN key[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 46.040000 248.850000 46.110000 248.920000 ;
    END
  END key[43]
  PIN key[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 45.090000 248.850000 45.160000 248.920000 ;
    END
  END key[42]
  PIN key[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 44.140000 248.850000 44.210000 248.920000 ;
    END
  END key[41]
  PIN key[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 43.190000 248.850000 43.260000 248.920000 ;
    END
  END key[40]
  PIN key[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 42.240000 248.850000 42.310000 248.920000 ;
    END
  END key[39]
  PIN key[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 41.290000 248.850000 41.360000 248.920000 ;
    END
  END key[38]
  PIN key[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 40.340000 248.850000 40.410000 248.920000 ;
    END
  END key[37]
  PIN key[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 39.390000 248.850000 39.460000 248.920000 ;
    END
  END key[36]
  PIN key[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 38.440000 248.850000 38.510000 248.920000 ;
    END
  END key[35]
  PIN key[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 37.490000 248.850000 37.560000 248.920000 ;
    END
  END key[34]
  PIN key[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 36.540000 248.850000 36.610000 248.920000 ;
    END
  END key[33]
  PIN key[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 35.590000 248.850000 35.660000 248.920000 ;
    END
  END key[32]
  PIN key[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 34.640000 248.850000 34.710000 248.920000 ;
    END
  END key[31]
  PIN key[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 33.690000 248.850000 33.760000 248.920000 ;
    END
  END key[30]
  PIN key[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 32.740000 248.850000 32.810000 248.920000 ;
    END
  END key[29]
  PIN key[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 31.790000 248.850000 31.860000 248.920000 ;
    END
  END key[28]
  PIN key[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 30.840000 248.850000 30.910000 248.920000 ;
    END
  END key[27]
  PIN key[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 29.890000 248.850000 29.960000 248.920000 ;
    END
  END key[26]
  PIN key[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 28.940000 248.850000 29.010000 248.920000 ;
    END
  END key[25]
  PIN key[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 27.990000 248.850000 28.060000 248.920000 ;
    END
  END key[24]
  PIN key[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 27.040000 248.850000 27.110000 248.920000 ;
    END
  END key[23]
  PIN key[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 26.090000 248.850000 26.160000 248.920000 ;
    END
  END key[22]
  PIN key[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 25.140000 248.850000 25.210000 248.920000 ;
    END
  END key[21]
  PIN key[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 24.190000 248.850000 24.260000 248.920000 ;
    END
  END key[20]
  PIN key[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 23.240000 248.850000 23.310000 248.920000 ;
    END
  END key[19]
  PIN key[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 22.290000 248.850000 22.360000 248.920000 ;
    END
  END key[18]
  PIN key[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 21.340000 248.850000 21.410000 248.920000 ;
    END
  END key[17]
  PIN key[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 20.390000 248.850000 20.460000 248.920000 ;
    END
  END key[16]
  PIN key[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 19.440000 248.850000 19.510000 248.920000 ;
    END
  END key[15]
  PIN key[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 18.490000 248.850000 18.560000 248.920000 ;
    END
  END key[14]
  PIN key[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 17.540000 248.850000 17.610000 248.920000 ;
    END
  END key[13]
  PIN key[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 16.590000 248.850000 16.660000 248.920000 ;
    END
  END key[12]
  PIN key[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 15.640000 248.850000 15.710000 248.920000 ;
    END
  END key[11]
  PIN key[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 14.690000 248.850000 14.760000 248.920000 ;
    END
  END key[10]
  PIN key[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 13.740000 248.850000 13.810000 248.920000 ;
    END
  END key[9]
  PIN key[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 12.790000 248.850000 12.860000 248.920000 ;
    END
  END key[8]
  PIN key[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 11.840000 248.850000 11.910000 248.920000 ;
    END
  END key[7]
  PIN key[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 10.890000 248.850000 10.960000 248.920000 ;
    END
  END key[6]
  PIN key[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.940000 248.850000 10.010000 248.920000 ;
    END
  END key[5]
  PIN key[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 8.990000 248.850000 9.060000 248.920000 ;
    END
  END key[4]
  PIN key[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 8.040000 248.850000 8.110000 248.920000 ;
    END
  END key[3]
  PIN key[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 7.090000 248.850000 7.160000 248.920000 ;
    END
  END key[2]
  PIN key[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 6.140000 248.850000 6.210000 248.920000 ;
    END
  END key[1]
  PIN key[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 5.190000 248.850000 5.260000 248.920000 ;
    END
  END key[0]
  PIN plain[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 247.440000 248.850000 247.510000 248.920000 ;
    END
  END plain[127]
  PIN plain[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 246.490000 248.850000 246.560000 248.920000 ;
    END
  END plain[126]
  PIN plain[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 245.540000 248.850000 245.610000 248.920000 ;
    END
  END plain[125]
  PIN plain[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 244.590000 248.850000 244.660000 248.920000 ;
    END
  END plain[124]
  PIN plain[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 243.640000 248.850000 243.710000 248.920000 ;
    END
  END plain[123]
  PIN plain[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 242.690000 248.850000 242.760000 248.920000 ;
    END
  END plain[122]
  PIN plain[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 241.740000 248.850000 241.810000 248.920000 ;
    END
  END plain[121]
  PIN plain[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 240.790000 248.850000 240.860000 248.920000 ;
    END
  END plain[120]
  PIN plain[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 239.840000 248.850000 239.910000 248.920000 ;
    END
  END plain[119]
  PIN plain[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 238.890000 248.850000 238.960000 248.920000 ;
    END
  END plain[118]
  PIN plain[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 237.940000 248.850000 238.010000 248.920000 ;
    END
  END plain[117]
  PIN plain[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 236.990000 248.850000 237.060000 248.920000 ;
    END
  END plain[116]
  PIN plain[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 236.040000 248.850000 236.110000 248.920000 ;
    END
  END plain[115]
  PIN plain[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 235.090000 248.850000 235.160000 248.920000 ;
    END
  END plain[114]
  PIN plain[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 234.140000 248.850000 234.210000 248.920000 ;
    END
  END plain[113]
  PIN plain[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 233.190000 248.850000 233.260000 248.920000 ;
    END
  END plain[112]
  PIN plain[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 232.240000 248.850000 232.310000 248.920000 ;
    END
  END plain[111]
  PIN plain[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 231.290000 248.850000 231.360000 248.920000 ;
    END
  END plain[110]
  PIN plain[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 230.340000 248.850000 230.410000 248.920000 ;
    END
  END plain[109]
  PIN plain[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 229.390000 248.850000 229.460000 248.920000 ;
    END
  END plain[108]
  PIN plain[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 228.440000 248.850000 228.510000 248.920000 ;
    END
  END plain[107]
  PIN plain[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 227.490000 248.850000 227.560000 248.920000 ;
    END
  END plain[106]
  PIN plain[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 226.540000 248.850000 226.610000 248.920000 ;
    END
  END plain[105]
  PIN plain[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 225.590000 248.850000 225.660000 248.920000 ;
    END
  END plain[104]
  PIN plain[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 224.640000 248.850000 224.710000 248.920000 ;
    END
  END plain[103]
  PIN plain[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 223.690000 248.850000 223.760000 248.920000 ;
    END
  END plain[102]
  PIN plain[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 222.740000 248.850000 222.810000 248.920000 ;
    END
  END plain[101]
  PIN plain[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 221.790000 248.850000 221.860000 248.920000 ;
    END
  END plain[100]
  PIN plain[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 220.840000 248.850000 220.910000 248.920000 ;
    END
  END plain[99]
  PIN plain[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 219.890000 248.850000 219.960000 248.920000 ;
    END
  END plain[98]
  PIN plain[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 218.940000 248.850000 219.010000 248.920000 ;
    END
  END plain[97]
  PIN plain[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 217.990000 248.850000 218.060000 248.920000 ;
    END
  END plain[96]
  PIN plain[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 217.040000 248.850000 217.110000 248.920000 ;
    END
  END plain[95]
  PIN plain[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 216.090000 248.850000 216.160000 248.920000 ;
    END
  END plain[94]
  PIN plain[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 215.140000 248.850000 215.210000 248.920000 ;
    END
  END plain[93]
  PIN plain[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 214.190000 248.850000 214.260000 248.920000 ;
    END
  END plain[92]
  PIN plain[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 213.240000 248.850000 213.310000 248.920000 ;
    END
  END plain[91]
  PIN plain[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 212.290000 248.850000 212.360000 248.920000 ;
    END
  END plain[90]
  PIN plain[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 211.340000 248.850000 211.410000 248.920000 ;
    END
  END plain[89]
  PIN plain[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 210.390000 248.850000 210.460000 248.920000 ;
    END
  END plain[88]
  PIN plain[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 209.440000 248.850000 209.510000 248.920000 ;
    END
  END plain[87]
  PIN plain[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 208.490000 248.850000 208.560000 248.920000 ;
    END
  END plain[86]
  PIN plain[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 207.540000 248.850000 207.610000 248.920000 ;
    END
  END plain[85]
  PIN plain[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 206.590000 248.850000 206.660000 248.920000 ;
    END
  END plain[84]
  PIN plain[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 205.640000 248.850000 205.710000 248.920000 ;
    END
  END plain[83]
  PIN plain[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 204.690000 248.850000 204.760000 248.920000 ;
    END
  END plain[82]
  PIN plain[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 203.740000 248.850000 203.810000 248.920000 ;
    END
  END plain[81]
  PIN plain[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 202.790000 248.850000 202.860000 248.920000 ;
    END
  END plain[80]
  PIN plain[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 201.840000 248.850000 201.910000 248.920000 ;
    END
  END plain[79]
  PIN plain[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 200.890000 248.850000 200.960000 248.920000 ;
    END
  END plain[78]
  PIN plain[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 199.940000 248.850000 200.010000 248.920000 ;
    END
  END plain[77]
  PIN plain[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 198.990000 248.850000 199.060000 248.920000 ;
    END
  END plain[76]
  PIN plain[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 198.040000 248.850000 198.110000 248.920000 ;
    END
  END plain[75]
  PIN plain[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 197.090000 248.850000 197.160000 248.920000 ;
    END
  END plain[74]
  PIN plain[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 196.140000 248.850000 196.210000 248.920000 ;
    END
  END plain[73]
  PIN plain[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 195.190000 248.850000 195.260000 248.920000 ;
    END
  END plain[72]
  PIN plain[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 194.240000 248.850000 194.310000 248.920000 ;
    END
  END plain[71]
  PIN plain[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 193.290000 248.850000 193.360000 248.920000 ;
    END
  END plain[70]
  PIN plain[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 192.340000 248.850000 192.410000 248.920000 ;
    END
  END plain[69]
  PIN plain[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 191.390000 248.850000 191.460000 248.920000 ;
    END
  END plain[68]
  PIN plain[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 190.440000 248.850000 190.510000 248.920000 ;
    END
  END plain[67]
  PIN plain[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 189.490000 248.850000 189.560000 248.920000 ;
    END
  END plain[66]
  PIN plain[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 188.540000 248.850000 188.610000 248.920000 ;
    END
  END plain[65]
  PIN plain[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 187.590000 248.850000 187.660000 248.920000 ;
    END
  END plain[64]
  PIN plain[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 186.640000 248.850000 186.710000 248.920000 ;
    END
  END plain[63]
  PIN plain[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 185.690000 248.850000 185.760000 248.920000 ;
    END
  END plain[62]
  PIN plain[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 184.740000 248.850000 184.810000 248.920000 ;
    END
  END plain[61]
  PIN plain[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 183.790000 248.850000 183.860000 248.920000 ;
    END
  END plain[60]
  PIN plain[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 182.840000 248.850000 182.910000 248.920000 ;
    END
  END plain[59]
  PIN plain[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 181.890000 248.850000 181.960000 248.920000 ;
    END
  END plain[58]
  PIN plain[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 180.940000 248.850000 181.010000 248.920000 ;
    END
  END plain[57]
  PIN plain[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 179.990000 248.850000 180.060000 248.920000 ;
    END
  END plain[56]
  PIN plain[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 179.040000 248.850000 179.110000 248.920000 ;
    END
  END plain[55]
  PIN plain[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 178.090000 248.850000 178.160000 248.920000 ;
    END
  END plain[54]
  PIN plain[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 177.140000 248.850000 177.210000 248.920000 ;
    END
  END plain[53]
  PIN plain[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 176.190000 248.850000 176.260000 248.920000 ;
    END
  END plain[52]
  PIN plain[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 175.240000 248.850000 175.310000 248.920000 ;
    END
  END plain[51]
  PIN plain[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 174.290000 248.850000 174.360000 248.920000 ;
    END
  END plain[50]
  PIN plain[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 173.340000 248.850000 173.410000 248.920000 ;
    END
  END plain[49]
  PIN plain[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 172.390000 248.850000 172.460000 248.920000 ;
    END
  END plain[48]
  PIN plain[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 171.440000 248.850000 171.510000 248.920000 ;
    END
  END plain[47]
  PIN plain[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 170.490000 248.850000 170.560000 248.920000 ;
    END
  END plain[46]
  PIN plain[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 169.540000 248.850000 169.610000 248.920000 ;
    END
  END plain[45]
  PIN plain[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.590000 248.850000 168.660000 248.920000 ;
    END
  END plain[44]
  PIN plain[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 167.640000 248.850000 167.710000 248.920000 ;
    END
  END plain[43]
  PIN plain[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 166.690000 248.850000 166.760000 248.920000 ;
    END
  END plain[42]
  PIN plain[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 165.740000 248.850000 165.810000 248.920000 ;
    END
  END plain[41]
  PIN plain[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 164.790000 248.850000 164.860000 248.920000 ;
    END
  END plain[40]
  PIN plain[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 163.840000 248.850000 163.910000 248.920000 ;
    END
  END plain[39]
  PIN plain[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 162.890000 248.850000 162.960000 248.920000 ;
    END
  END plain[38]
  PIN plain[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 161.940000 248.850000 162.010000 248.920000 ;
    END
  END plain[37]
  PIN plain[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 160.990000 248.850000 161.060000 248.920000 ;
    END
  END plain[36]
  PIN plain[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 160.040000 248.850000 160.110000 248.920000 ;
    END
  END plain[35]
  PIN plain[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 159.090000 248.850000 159.160000 248.920000 ;
    END
  END plain[34]
  PIN plain[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 158.140000 248.850000 158.210000 248.920000 ;
    END
  END plain[33]
  PIN plain[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 157.190000 248.850000 157.260000 248.920000 ;
    END
  END plain[32]
  PIN plain[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 156.240000 248.850000 156.310000 248.920000 ;
    END
  END plain[31]
  PIN plain[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 155.290000 248.850000 155.360000 248.920000 ;
    END
  END plain[30]
  PIN plain[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 154.340000 248.850000 154.410000 248.920000 ;
    END
  END plain[29]
  PIN plain[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 153.390000 248.850000 153.460000 248.920000 ;
    END
  END plain[28]
  PIN plain[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 152.440000 248.850000 152.510000 248.920000 ;
    END
  END plain[27]
  PIN plain[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 151.490000 248.850000 151.560000 248.920000 ;
    END
  END plain[26]
  PIN plain[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 150.540000 248.850000 150.610000 248.920000 ;
    END
  END plain[25]
  PIN plain[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 149.590000 248.850000 149.660000 248.920000 ;
    END
  END plain[24]
  PIN plain[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 148.640000 248.850000 148.710000 248.920000 ;
    END
  END plain[23]
  PIN plain[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 147.690000 248.850000 147.760000 248.920000 ;
    END
  END plain[22]
  PIN plain[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 146.740000 248.850000 146.810000 248.920000 ;
    END
  END plain[21]
  PIN plain[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 145.790000 248.850000 145.860000 248.920000 ;
    END
  END plain[20]
  PIN plain[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 144.840000 248.850000 144.910000 248.920000 ;
    END
  END plain[19]
  PIN plain[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 143.890000 248.850000 143.960000 248.920000 ;
    END
  END plain[18]
  PIN plain[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 142.940000 248.850000 143.010000 248.920000 ;
    END
  END plain[17]
  PIN plain[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 141.990000 248.850000 142.060000 248.920000 ;
    END
  END plain[16]
  PIN plain[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 141.040000 248.850000 141.110000 248.920000 ;
    END
  END plain[15]
  PIN plain[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 140.090000 248.850000 140.160000 248.920000 ;
    END
  END plain[14]
  PIN plain[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 139.140000 248.850000 139.210000 248.920000 ;
    END
  END plain[13]
  PIN plain[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 138.190000 248.850000 138.260000 248.920000 ;
    END
  END plain[12]
  PIN plain[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 137.240000 248.850000 137.310000 248.920000 ;
    END
  END plain[11]
  PIN plain[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 136.290000 248.850000 136.360000 248.920000 ;
    END
  END plain[10]
  PIN plain[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 135.340000 248.850000 135.410000 248.920000 ;
    END
  END plain[9]
  PIN plain[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 134.390000 248.850000 134.460000 248.920000 ;
    END
  END plain[8]
  PIN plain[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 133.440000 248.850000 133.510000 248.920000 ;
    END
  END plain[7]
  PIN plain[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 132.490000 248.850000 132.560000 248.920000 ;
    END
  END plain[6]
  PIN plain[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 131.540000 248.850000 131.610000 248.920000 ;
    END
  END plain[5]
  PIN plain[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 130.590000 248.850000 130.660000 248.920000 ;
    END
  END plain[4]
  PIN plain[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 129.640000 248.850000 129.710000 248.920000 ;
    END
  END plain[3]
  PIN plain[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 128.690000 248.850000 128.760000 248.920000 ;
    END
  END plain[2]
  PIN plain[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 127.740000 248.850000 127.810000 248.920000 ;
    END
  END plain[1]
  PIN plain[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 126.790000 248.850000 126.860000 248.920000 ;
    END
  END plain[0]
  PIN ready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 246.300000 0.000000 246.370000 0.070000 ;
    END
  END ready
  PIN cipher[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.100000 0.000000 3.170000 0.070000 ;
    END
  END cipher[127]
  PIN cipher[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 5.000000 0.000000 5.070000 0.070000 ;
    END
  END cipher[126]
  PIN cipher[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 6.900000 0.000000 6.970000 0.070000 ;
    END
  END cipher[125]
  PIN cipher[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 8.800000 0.000000 8.870000 0.070000 ;
    END
  END cipher[124]
  PIN cipher[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 10.700000 0.000000 10.770000 0.070000 ;
    END
  END cipher[123]
  PIN cipher[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 12.600000 0.000000 12.670000 0.070000 ;
    END
  END cipher[122]
  PIN cipher[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 14.500000 0.000000 14.570000 0.070000 ;
    END
  END cipher[121]
  PIN cipher[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 16.400000 0.000000 16.470000 0.070000 ;
    END
  END cipher[120]
  PIN cipher[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 18.300000 0.000000 18.370000 0.070000 ;
    END
  END cipher[119]
  PIN cipher[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 20.200000 0.000000 20.270000 0.070000 ;
    END
  END cipher[118]
  PIN cipher[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 22.100000 0.000000 22.170000 0.070000 ;
    END
  END cipher[117]
  PIN cipher[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 24.000000 0.000000 24.070000 0.070000 ;
    END
  END cipher[116]
  PIN cipher[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 25.900000 0.000000 25.970000 0.070000 ;
    END
  END cipher[115]
  PIN cipher[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 27.800000 0.000000 27.870000 0.070000 ;
    END
  END cipher[114]
  PIN cipher[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 29.700000 0.000000 29.770000 0.070000 ;
    END
  END cipher[113]
  PIN cipher[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 31.600000 0.000000 31.670000 0.070000 ;
    END
  END cipher[112]
  PIN cipher[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 33.500000 0.000000 33.570000 0.070000 ;
    END
  END cipher[111]
  PIN cipher[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 35.400000 0.000000 35.470000 0.070000 ;
    END
  END cipher[110]
  PIN cipher[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 37.300000 0.000000 37.370000 0.070000 ;
    END
  END cipher[109]
  PIN cipher[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 39.200000 0.000000 39.270000 0.070000 ;
    END
  END cipher[108]
  PIN cipher[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 41.100000 0.000000 41.170000 0.070000 ;
    END
  END cipher[107]
  PIN cipher[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 43.000000 0.000000 43.070000 0.070000 ;
    END
  END cipher[106]
  PIN cipher[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 44.900000 0.000000 44.970000 0.070000 ;
    END
  END cipher[105]
  PIN cipher[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 46.800000 0.000000 46.870000 0.070000 ;
    END
  END cipher[104]
  PIN cipher[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 48.700000 0.000000 48.770000 0.070000 ;
    END
  END cipher[103]
  PIN cipher[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 50.600000 0.000000 50.670000 0.070000 ;
    END
  END cipher[102]
  PIN cipher[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 52.500000 0.000000 52.570000 0.070000 ;
    END
  END cipher[101]
  PIN cipher[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 54.400000 0.000000 54.470000 0.070000 ;
    END
  END cipher[100]
  PIN cipher[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 56.300000 0.000000 56.370000 0.070000 ;
    END
  END cipher[99]
  PIN cipher[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 58.200000 0.000000 58.270000 0.070000 ;
    END
  END cipher[98]
  PIN cipher[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 60.100000 0.000000 60.170000 0.070000 ;
    END
  END cipher[97]
  PIN cipher[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 62.000000 0.000000 62.070000 0.070000 ;
    END
  END cipher[96]
  PIN cipher[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 63.900000 0.000000 63.970000 0.070000 ;
    END
  END cipher[95]
  PIN cipher[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 65.800000 0.000000 65.870000 0.070000 ;
    END
  END cipher[94]
  PIN cipher[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 67.700000 0.000000 67.770000 0.070000 ;
    END
  END cipher[93]
  PIN cipher[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 69.600000 0.000000 69.670000 0.070000 ;
    END
  END cipher[92]
  PIN cipher[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 71.500000 0.000000 71.570000 0.070000 ;
    END
  END cipher[91]
  PIN cipher[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 73.400000 0.000000 73.470000 0.070000 ;
    END
  END cipher[90]
  PIN cipher[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 75.300000 0.000000 75.370000 0.070000 ;
    END
  END cipher[89]
  PIN cipher[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 77.200000 0.000000 77.270000 0.070000 ;
    END
  END cipher[88]
  PIN cipher[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 79.100000 0.000000 79.170000 0.070000 ;
    END
  END cipher[87]
  PIN cipher[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 81.000000 0.000000 81.070000 0.070000 ;
    END
  END cipher[86]
  PIN cipher[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 82.900000 0.000000 82.970000 0.070000 ;
    END
  END cipher[85]
  PIN cipher[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 84.800000 0.000000 84.870000 0.070000 ;
    END
  END cipher[84]
  PIN cipher[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 86.700000 0.000000 86.770000 0.070000 ;
    END
  END cipher[83]
  PIN cipher[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 88.600000 0.000000 88.670000 0.070000 ;
    END
  END cipher[82]
  PIN cipher[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 90.500000 0.000000 90.570000 0.070000 ;
    END
  END cipher[81]
  PIN cipher[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 92.400000 0.000000 92.470000 0.070000 ;
    END
  END cipher[80]
  PIN cipher[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 94.300000 0.000000 94.370000 0.070000 ;
    END
  END cipher[79]
  PIN cipher[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 96.200000 0.000000 96.270000 0.070000 ;
    END
  END cipher[78]
  PIN cipher[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 98.100000 0.000000 98.170000 0.070000 ;
    END
  END cipher[77]
  PIN cipher[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 100.000000 0.000000 100.070000 0.070000 ;
    END
  END cipher[76]
  PIN cipher[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 101.900000 0.000000 101.970000 0.070000 ;
    END
  END cipher[75]
  PIN cipher[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 103.800000 0.000000 103.870000 0.070000 ;
    END
  END cipher[74]
  PIN cipher[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 105.700000 0.000000 105.770000 0.070000 ;
    END
  END cipher[73]
  PIN cipher[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 107.600000 0.000000 107.670000 0.070000 ;
    END
  END cipher[72]
  PIN cipher[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 109.500000 0.000000 109.570000 0.070000 ;
    END
  END cipher[71]
  PIN cipher[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 111.400000 0.000000 111.470000 0.070000 ;
    END
  END cipher[70]
  PIN cipher[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 113.300000 0.000000 113.370000 0.070000 ;
    END
  END cipher[69]
  PIN cipher[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 115.200000 0.000000 115.270000 0.070000 ;
    END
  END cipher[68]
  PIN cipher[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 117.100000 0.000000 117.170000 0.070000 ;
    END
  END cipher[67]
  PIN cipher[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 119.000000 0.000000 119.070000 0.070000 ;
    END
  END cipher[66]
  PIN cipher[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 120.900000 0.000000 120.970000 0.070000 ;
    END
  END cipher[65]
  PIN cipher[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 122.800000 0.000000 122.870000 0.070000 ;
    END
  END cipher[64]
  PIN cipher[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 124.700000 0.000000 124.770000 0.070000 ;
    END
  END cipher[63]
  PIN cipher[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 126.600000 0.000000 126.670000 0.070000 ;
    END
  END cipher[62]
  PIN cipher[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 128.500000 0.000000 128.570000 0.070000 ;
    END
  END cipher[61]
  PIN cipher[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 130.400000 0.000000 130.470000 0.070000 ;
    END
  END cipher[60]
  PIN cipher[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 132.300000 0.000000 132.370000 0.070000 ;
    END
  END cipher[59]
  PIN cipher[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 134.200000 0.000000 134.270000 0.070000 ;
    END
  END cipher[58]
  PIN cipher[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 136.100000 0.000000 136.170000 0.070000 ;
    END
  END cipher[57]
  PIN cipher[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 138.000000 0.000000 138.070000 0.070000 ;
    END
  END cipher[56]
  PIN cipher[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 139.900000 0.000000 139.970000 0.070000 ;
    END
  END cipher[55]
  PIN cipher[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 141.800000 0.000000 141.870000 0.070000 ;
    END
  END cipher[54]
  PIN cipher[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 143.700000 0.000000 143.770000 0.070000 ;
    END
  END cipher[53]
  PIN cipher[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 145.600000 0.000000 145.670000 0.070000 ;
    END
  END cipher[52]
  PIN cipher[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 147.500000 0.000000 147.570000 0.070000 ;
    END
  END cipher[51]
  PIN cipher[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 149.400000 0.000000 149.470000 0.070000 ;
    END
  END cipher[50]
  PIN cipher[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 151.300000 0.000000 151.370000 0.070000 ;
    END
  END cipher[49]
  PIN cipher[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 153.200000 0.000000 153.270000 0.070000 ;
    END
  END cipher[48]
  PIN cipher[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 155.100000 0.000000 155.170000 0.070000 ;
    END
  END cipher[47]
  PIN cipher[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 157.000000 0.000000 157.070000 0.070000 ;
    END
  END cipher[46]
  PIN cipher[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 158.900000 0.000000 158.970000 0.070000 ;
    END
  END cipher[45]
  PIN cipher[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 160.800000 0.000000 160.870000 0.070000 ;
    END
  END cipher[44]
  PIN cipher[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 162.700000 0.000000 162.770000 0.070000 ;
    END
  END cipher[43]
  PIN cipher[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 164.600000 0.000000 164.670000 0.070000 ;
    END
  END cipher[42]
  PIN cipher[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 166.500000 0.000000 166.570000 0.070000 ;
    END
  END cipher[41]
  PIN cipher[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.400000 0.000000 168.470000 0.070000 ;
    END
  END cipher[40]
  PIN cipher[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 170.300000 0.000000 170.370000 0.070000 ;
    END
  END cipher[39]
  PIN cipher[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 172.200000 0.000000 172.270000 0.070000 ;
    END
  END cipher[38]
  PIN cipher[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 174.100000 0.000000 174.170000 0.070000 ;
    END
  END cipher[37]
  PIN cipher[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 176.000000 0.000000 176.070000 0.070000 ;
    END
  END cipher[36]
  PIN cipher[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 177.900000 0.000000 177.970000 0.070000 ;
    END
  END cipher[35]
  PIN cipher[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 179.800000 0.000000 179.870000 0.070000 ;
    END
  END cipher[34]
  PIN cipher[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 181.700000 0.000000 181.770000 0.070000 ;
    END
  END cipher[33]
  PIN cipher[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 183.600000 0.000000 183.670000 0.070000 ;
    END
  END cipher[32]
  PIN cipher[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 185.500000 0.000000 185.570000 0.070000 ;
    END
  END cipher[31]
  PIN cipher[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 187.400000 0.000000 187.470000 0.070000 ;
    END
  END cipher[30]
  PIN cipher[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 189.300000 0.000000 189.370000 0.070000 ;
    END
  END cipher[29]
  PIN cipher[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 191.200000 0.000000 191.270000 0.070000 ;
    END
  END cipher[28]
  PIN cipher[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 193.100000 0.000000 193.170000 0.070000 ;
    END
  END cipher[27]
  PIN cipher[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 195.000000 0.000000 195.070000 0.070000 ;
    END
  END cipher[26]
  PIN cipher[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 196.900000 0.000000 196.970000 0.070000 ;
    END
  END cipher[25]
  PIN cipher[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 198.800000 0.000000 198.870000 0.070000 ;
    END
  END cipher[24]
  PIN cipher[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 200.700000 0.000000 200.770000 0.070000 ;
    END
  END cipher[23]
  PIN cipher[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 202.600000 0.000000 202.670000 0.070000 ;
    END
  END cipher[22]
  PIN cipher[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 204.500000 0.000000 204.570000 0.070000 ;
    END
  END cipher[21]
  PIN cipher[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 206.400000 0.000000 206.470000 0.070000 ;
    END
  END cipher[20]
  PIN cipher[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 208.300000 0.000000 208.370000 0.070000 ;
    END
  END cipher[19]
  PIN cipher[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 210.200000 0.000000 210.270000 0.070000 ;
    END
  END cipher[18]
  PIN cipher[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 212.100000 0.000000 212.170000 0.070000 ;
    END
  END cipher[17]
  PIN cipher[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 214.000000 0.000000 214.070000 0.070000 ;
    END
  END cipher[16]
  PIN cipher[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 215.900000 0.000000 215.970000 0.070000 ;
    END
  END cipher[15]
  PIN cipher[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 217.800000 0.000000 217.870000 0.070000 ;
    END
  END cipher[14]
  PIN cipher[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 219.700000 0.000000 219.770000 0.070000 ;
    END
  END cipher[13]
  PIN cipher[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 221.600000 0.000000 221.670000 0.070000 ;
    END
  END cipher[12]
  PIN cipher[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 223.500000 0.000000 223.570000 0.070000 ;
    END
  END cipher[11]
  PIN cipher[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 225.400000 0.000000 225.470000 0.070000 ;
    END
  END cipher[10]
  PIN cipher[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 227.300000 0.000000 227.370000 0.070000 ;
    END
  END cipher[9]
  PIN cipher[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 229.200000 0.000000 229.270000 0.070000 ;
    END
  END cipher[8]
  PIN cipher[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 231.100000 0.000000 231.170000 0.070000 ;
    END
  END cipher[7]
  PIN cipher[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 233.000000 0.000000 233.070000 0.070000 ;
    END
  END cipher[6]
  PIN cipher[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 234.900000 0.000000 234.970000 0.070000 ;
    END
  END cipher[5]
  PIN cipher[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 236.800000 0.000000 236.870000 0.070000 ;
    END
  END cipher[4]
  PIN cipher[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 238.700000 0.000000 238.770000 0.070000 ;
    END
  END cipher[3]
  PIN cipher[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 240.600000 0.000000 240.670000 0.070000 ;
    END
  END cipher[2]
  PIN cipher[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 242.500000 0.000000 242.570000 0.070000 ;
    END
  END cipher[1]
  PIN cipher[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 244.400000 0.000000 244.470000 0.070000 ;
    END
  END cipher[0]
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 251.180000 248.920000 ;
    LAYER metal2 ;
      RECT 247.580000 248.780000 251.180000 248.920000 ;
      RECT 246.630000 248.780000 247.370000 248.920000 ;
      RECT 245.680000 248.780000 246.420000 248.920000 ;
      RECT 244.730000 248.780000 245.470000 248.920000 ;
      RECT 243.780000 248.780000 244.520000 248.920000 ;
      RECT 242.830000 248.780000 243.570000 248.920000 ;
      RECT 241.880000 248.780000 242.620000 248.920000 ;
      RECT 240.930000 248.780000 241.670000 248.920000 ;
      RECT 239.980000 248.780000 240.720000 248.920000 ;
      RECT 239.030000 248.780000 239.770000 248.920000 ;
      RECT 238.080000 248.780000 238.820000 248.920000 ;
      RECT 237.130000 248.780000 237.870000 248.920000 ;
      RECT 236.180000 248.780000 236.920000 248.920000 ;
      RECT 235.230000 248.780000 235.970000 248.920000 ;
      RECT 234.280000 248.780000 235.020000 248.920000 ;
      RECT 233.330000 248.780000 234.070000 248.920000 ;
      RECT 232.380000 248.780000 233.120000 248.920000 ;
      RECT 231.430000 248.780000 232.170000 248.920000 ;
      RECT 230.480000 248.780000 231.220000 248.920000 ;
      RECT 229.530000 248.780000 230.270000 248.920000 ;
      RECT 228.580000 248.780000 229.320000 248.920000 ;
      RECT 227.630000 248.780000 228.370000 248.920000 ;
      RECT 226.680000 248.780000 227.420000 248.920000 ;
      RECT 225.730000 248.780000 226.470000 248.920000 ;
      RECT 224.780000 248.780000 225.520000 248.920000 ;
      RECT 223.830000 248.780000 224.570000 248.920000 ;
      RECT 222.880000 248.780000 223.620000 248.920000 ;
      RECT 221.930000 248.780000 222.670000 248.920000 ;
      RECT 220.980000 248.780000 221.720000 248.920000 ;
      RECT 220.030000 248.780000 220.770000 248.920000 ;
      RECT 219.080000 248.780000 219.820000 248.920000 ;
      RECT 218.130000 248.780000 218.870000 248.920000 ;
      RECT 217.180000 248.780000 217.920000 248.920000 ;
      RECT 216.230000 248.780000 216.970000 248.920000 ;
      RECT 215.280000 248.780000 216.020000 248.920000 ;
      RECT 214.330000 248.780000 215.070000 248.920000 ;
      RECT 213.380000 248.780000 214.120000 248.920000 ;
      RECT 212.430000 248.780000 213.170000 248.920000 ;
      RECT 211.480000 248.780000 212.220000 248.920000 ;
      RECT 210.530000 248.780000 211.270000 248.920000 ;
      RECT 209.580000 248.780000 210.320000 248.920000 ;
      RECT 208.630000 248.780000 209.370000 248.920000 ;
      RECT 207.680000 248.780000 208.420000 248.920000 ;
      RECT 206.730000 248.780000 207.470000 248.920000 ;
      RECT 205.780000 248.780000 206.520000 248.920000 ;
      RECT 204.830000 248.780000 205.570000 248.920000 ;
      RECT 203.880000 248.780000 204.620000 248.920000 ;
      RECT 202.930000 248.780000 203.670000 248.920000 ;
      RECT 201.980000 248.780000 202.720000 248.920000 ;
      RECT 201.030000 248.780000 201.770000 248.920000 ;
      RECT 200.080000 248.780000 200.820000 248.920000 ;
      RECT 199.130000 248.780000 199.870000 248.920000 ;
      RECT 198.180000 248.780000 198.920000 248.920000 ;
      RECT 197.230000 248.780000 197.970000 248.920000 ;
      RECT 196.280000 248.780000 197.020000 248.920000 ;
      RECT 195.330000 248.780000 196.070000 248.920000 ;
      RECT 194.380000 248.780000 195.120000 248.920000 ;
      RECT 193.430000 248.780000 194.170000 248.920000 ;
      RECT 192.480000 248.780000 193.220000 248.920000 ;
      RECT 191.530000 248.780000 192.270000 248.920000 ;
      RECT 190.580000 248.780000 191.320000 248.920000 ;
      RECT 189.630000 248.780000 190.370000 248.920000 ;
      RECT 188.680000 248.780000 189.420000 248.920000 ;
      RECT 187.730000 248.780000 188.470000 248.920000 ;
      RECT 186.780000 248.780000 187.520000 248.920000 ;
      RECT 185.830000 248.780000 186.570000 248.920000 ;
      RECT 184.880000 248.780000 185.620000 248.920000 ;
      RECT 183.930000 248.780000 184.670000 248.920000 ;
      RECT 182.980000 248.780000 183.720000 248.920000 ;
      RECT 182.030000 248.780000 182.770000 248.920000 ;
      RECT 181.080000 248.780000 181.820000 248.920000 ;
      RECT 180.130000 248.780000 180.870000 248.920000 ;
      RECT 179.180000 248.780000 179.920000 248.920000 ;
      RECT 178.230000 248.780000 178.970000 248.920000 ;
      RECT 177.280000 248.780000 178.020000 248.920000 ;
      RECT 176.330000 248.780000 177.070000 248.920000 ;
      RECT 175.380000 248.780000 176.120000 248.920000 ;
      RECT 174.430000 248.780000 175.170000 248.920000 ;
      RECT 173.480000 248.780000 174.220000 248.920000 ;
      RECT 172.530000 248.780000 173.270000 248.920000 ;
      RECT 171.580000 248.780000 172.320000 248.920000 ;
      RECT 170.630000 248.780000 171.370000 248.920000 ;
      RECT 169.680000 248.780000 170.420000 248.920000 ;
      RECT 168.730000 248.780000 169.470000 248.920000 ;
      RECT 167.780000 248.780000 168.520000 248.920000 ;
      RECT 166.830000 248.780000 167.570000 248.920000 ;
      RECT 165.880000 248.780000 166.620000 248.920000 ;
      RECT 164.930000 248.780000 165.670000 248.920000 ;
      RECT 163.980000 248.780000 164.720000 248.920000 ;
      RECT 163.030000 248.780000 163.770000 248.920000 ;
      RECT 162.080000 248.780000 162.820000 248.920000 ;
      RECT 161.130000 248.780000 161.870000 248.920000 ;
      RECT 160.180000 248.780000 160.920000 248.920000 ;
      RECT 159.230000 248.780000 159.970000 248.920000 ;
      RECT 158.280000 248.780000 159.020000 248.920000 ;
      RECT 157.330000 248.780000 158.070000 248.920000 ;
      RECT 156.380000 248.780000 157.120000 248.920000 ;
      RECT 155.430000 248.780000 156.170000 248.920000 ;
      RECT 154.480000 248.780000 155.220000 248.920000 ;
      RECT 153.530000 248.780000 154.270000 248.920000 ;
      RECT 152.580000 248.780000 153.320000 248.920000 ;
      RECT 151.630000 248.780000 152.370000 248.920000 ;
      RECT 150.680000 248.780000 151.420000 248.920000 ;
      RECT 149.730000 248.780000 150.470000 248.920000 ;
      RECT 148.780000 248.780000 149.520000 248.920000 ;
      RECT 147.830000 248.780000 148.570000 248.920000 ;
      RECT 146.880000 248.780000 147.620000 248.920000 ;
      RECT 145.930000 248.780000 146.670000 248.920000 ;
      RECT 144.980000 248.780000 145.720000 248.920000 ;
      RECT 144.030000 248.780000 144.770000 248.920000 ;
      RECT 143.080000 248.780000 143.820000 248.920000 ;
      RECT 142.130000 248.780000 142.870000 248.920000 ;
      RECT 141.180000 248.780000 141.920000 248.920000 ;
      RECT 140.230000 248.780000 140.970000 248.920000 ;
      RECT 139.280000 248.780000 140.020000 248.920000 ;
      RECT 138.330000 248.780000 139.070000 248.920000 ;
      RECT 137.380000 248.780000 138.120000 248.920000 ;
      RECT 136.430000 248.780000 137.170000 248.920000 ;
      RECT 135.480000 248.780000 136.220000 248.920000 ;
      RECT 134.530000 248.780000 135.270000 248.920000 ;
      RECT 133.580000 248.780000 134.320000 248.920000 ;
      RECT 132.630000 248.780000 133.370000 248.920000 ;
      RECT 131.680000 248.780000 132.420000 248.920000 ;
      RECT 130.730000 248.780000 131.470000 248.920000 ;
      RECT 129.780000 248.780000 130.520000 248.920000 ;
      RECT 128.830000 248.780000 129.570000 248.920000 ;
      RECT 127.880000 248.780000 128.620000 248.920000 ;
      RECT 126.930000 248.780000 127.670000 248.920000 ;
      RECT 125.980000 248.780000 126.720000 248.920000 ;
      RECT 125.030000 248.780000 125.770000 248.920000 ;
      RECT 124.080000 248.780000 124.820000 248.920000 ;
      RECT 123.130000 248.780000 123.870000 248.920000 ;
      RECT 122.180000 248.780000 122.920000 248.920000 ;
      RECT 121.230000 248.780000 121.970000 248.920000 ;
      RECT 120.280000 248.780000 121.020000 248.920000 ;
      RECT 119.330000 248.780000 120.070000 248.920000 ;
      RECT 118.380000 248.780000 119.120000 248.920000 ;
      RECT 117.430000 248.780000 118.170000 248.920000 ;
      RECT 116.480000 248.780000 117.220000 248.920000 ;
      RECT 115.530000 248.780000 116.270000 248.920000 ;
      RECT 114.580000 248.780000 115.320000 248.920000 ;
      RECT 113.630000 248.780000 114.370000 248.920000 ;
      RECT 112.680000 248.780000 113.420000 248.920000 ;
      RECT 111.730000 248.780000 112.470000 248.920000 ;
      RECT 110.780000 248.780000 111.520000 248.920000 ;
      RECT 109.830000 248.780000 110.570000 248.920000 ;
      RECT 108.880000 248.780000 109.620000 248.920000 ;
      RECT 107.930000 248.780000 108.670000 248.920000 ;
      RECT 106.980000 248.780000 107.720000 248.920000 ;
      RECT 106.030000 248.780000 106.770000 248.920000 ;
      RECT 105.080000 248.780000 105.820000 248.920000 ;
      RECT 104.130000 248.780000 104.870000 248.920000 ;
      RECT 103.180000 248.780000 103.920000 248.920000 ;
      RECT 102.230000 248.780000 102.970000 248.920000 ;
      RECT 101.280000 248.780000 102.020000 248.920000 ;
      RECT 100.330000 248.780000 101.070000 248.920000 ;
      RECT 99.380000 248.780000 100.120000 248.920000 ;
      RECT 98.430000 248.780000 99.170000 248.920000 ;
      RECT 97.480000 248.780000 98.220000 248.920000 ;
      RECT 96.530000 248.780000 97.270000 248.920000 ;
      RECT 95.580000 248.780000 96.320000 248.920000 ;
      RECT 94.630000 248.780000 95.370000 248.920000 ;
      RECT 93.680000 248.780000 94.420000 248.920000 ;
      RECT 92.730000 248.780000 93.470000 248.920000 ;
      RECT 91.780000 248.780000 92.520000 248.920000 ;
      RECT 90.830000 248.780000 91.570000 248.920000 ;
      RECT 89.880000 248.780000 90.620000 248.920000 ;
      RECT 88.930000 248.780000 89.670000 248.920000 ;
      RECT 87.980000 248.780000 88.720000 248.920000 ;
      RECT 87.030000 248.780000 87.770000 248.920000 ;
      RECT 86.080000 248.780000 86.820000 248.920000 ;
      RECT 85.130000 248.780000 85.870000 248.920000 ;
      RECT 84.180000 248.780000 84.920000 248.920000 ;
      RECT 83.230000 248.780000 83.970000 248.920000 ;
      RECT 82.280000 248.780000 83.020000 248.920000 ;
      RECT 81.330000 248.780000 82.070000 248.920000 ;
      RECT 80.380000 248.780000 81.120000 248.920000 ;
      RECT 79.430000 248.780000 80.170000 248.920000 ;
      RECT 78.480000 248.780000 79.220000 248.920000 ;
      RECT 77.530000 248.780000 78.270000 248.920000 ;
      RECT 76.580000 248.780000 77.320000 248.920000 ;
      RECT 75.630000 248.780000 76.370000 248.920000 ;
      RECT 74.680000 248.780000 75.420000 248.920000 ;
      RECT 73.730000 248.780000 74.470000 248.920000 ;
      RECT 72.780000 248.780000 73.520000 248.920000 ;
      RECT 71.830000 248.780000 72.570000 248.920000 ;
      RECT 70.880000 248.780000 71.620000 248.920000 ;
      RECT 69.930000 248.780000 70.670000 248.920000 ;
      RECT 68.980000 248.780000 69.720000 248.920000 ;
      RECT 68.030000 248.780000 68.770000 248.920000 ;
      RECT 67.080000 248.780000 67.820000 248.920000 ;
      RECT 66.130000 248.780000 66.870000 248.920000 ;
      RECT 65.180000 248.780000 65.920000 248.920000 ;
      RECT 64.230000 248.780000 64.970000 248.920000 ;
      RECT 63.280000 248.780000 64.020000 248.920000 ;
      RECT 62.330000 248.780000 63.070000 248.920000 ;
      RECT 61.380000 248.780000 62.120000 248.920000 ;
      RECT 60.430000 248.780000 61.170000 248.920000 ;
      RECT 59.480000 248.780000 60.220000 248.920000 ;
      RECT 58.530000 248.780000 59.270000 248.920000 ;
      RECT 57.580000 248.780000 58.320000 248.920000 ;
      RECT 56.630000 248.780000 57.370000 248.920000 ;
      RECT 55.680000 248.780000 56.420000 248.920000 ;
      RECT 54.730000 248.780000 55.470000 248.920000 ;
      RECT 53.780000 248.780000 54.520000 248.920000 ;
      RECT 52.830000 248.780000 53.570000 248.920000 ;
      RECT 51.880000 248.780000 52.620000 248.920000 ;
      RECT 50.930000 248.780000 51.670000 248.920000 ;
      RECT 49.980000 248.780000 50.720000 248.920000 ;
      RECT 49.030000 248.780000 49.770000 248.920000 ;
      RECT 48.080000 248.780000 48.820000 248.920000 ;
      RECT 47.130000 248.780000 47.870000 248.920000 ;
      RECT 46.180000 248.780000 46.920000 248.920000 ;
      RECT 45.230000 248.780000 45.970000 248.920000 ;
      RECT 44.280000 248.780000 45.020000 248.920000 ;
      RECT 43.330000 248.780000 44.070000 248.920000 ;
      RECT 42.380000 248.780000 43.120000 248.920000 ;
      RECT 41.430000 248.780000 42.170000 248.920000 ;
      RECT 40.480000 248.780000 41.220000 248.920000 ;
      RECT 39.530000 248.780000 40.270000 248.920000 ;
      RECT 38.580000 248.780000 39.320000 248.920000 ;
      RECT 37.630000 248.780000 38.370000 248.920000 ;
      RECT 36.680000 248.780000 37.420000 248.920000 ;
      RECT 35.730000 248.780000 36.470000 248.920000 ;
      RECT 34.780000 248.780000 35.520000 248.920000 ;
      RECT 33.830000 248.780000 34.570000 248.920000 ;
      RECT 32.880000 248.780000 33.620000 248.920000 ;
      RECT 31.930000 248.780000 32.670000 248.920000 ;
      RECT 30.980000 248.780000 31.720000 248.920000 ;
      RECT 30.030000 248.780000 30.770000 248.920000 ;
      RECT 29.080000 248.780000 29.820000 248.920000 ;
      RECT 28.130000 248.780000 28.870000 248.920000 ;
      RECT 27.180000 248.780000 27.920000 248.920000 ;
      RECT 26.230000 248.780000 26.970000 248.920000 ;
      RECT 25.280000 248.780000 26.020000 248.920000 ;
      RECT 24.330000 248.780000 25.070000 248.920000 ;
      RECT 23.380000 248.780000 24.120000 248.920000 ;
      RECT 22.430000 248.780000 23.170000 248.920000 ;
      RECT 21.480000 248.780000 22.220000 248.920000 ;
      RECT 20.530000 248.780000 21.270000 248.920000 ;
      RECT 19.580000 248.780000 20.320000 248.920000 ;
      RECT 18.630000 248.780000 19.370000 248.920000 ;
      RECT 17.680000 248.780000 18.420000 248.920000 ;
      RECT 16.730000 248.780000 17.470000 248.920000 ;
      RECT 15.780000 248.780000 16.520000 248.920000 ;
      RECT 14.830000 248.780000 15.570000 248.920000 ;
      RECT 13.880000 248.780000 14.620000 248.920000 ;
      RECT 12.930000 248.780000 13.670000 248.920000 ;
      RECT 11.980000 248.780000 12.720000 248.920000 ;
      RECT 11.030000 248.780000 11.770000 248.920000 ;
      RECT 10.080000 248.780000 10.820000 248.920000 ;
      RECT 9.130000 248.780000 9.870000 248.920000 ;
      RECT 8.180000 248.780000 8.920000 248.920000 ;
      RECT 7.230000 248.780000 7.970000 248.920000 ;
      RECT 6.280000 248.780000 7.020000 248.920000 ;
      RECT 5.330000 248.780000 6.070000 248.920000 ;
      RECT 4.380000 248.780000 5.120000 248.920000 ;
      RECT 3.430000 248.780000 4.170000 248.920000 ;
      RECT 0.000000 248.780000 3.220000 248.920000 ;
      RECT 0.000000 0.140000 251.180000 248.780000 ;
      RECT 248.340000 0.000000 251.180000 0.140000 ;
      RECT 246.440000 0.000000 248.130000 0.140000 ;
      RECT 244.540000 0.000000 246.230000 0.140000 ;
      RECT 242.640000 0.000000 244.330000 0.140000 ;
      RECT 240.740000 0.000000 242.430000 0.140000 ;
      RECT 238.840000 0.000000 240.530000 0.140000 ;
      RECT 236.940000 0.000000 238.630000 0.140000 ;
      RECT 235.040000 0.000000 236.730000 0.140000 ;
      RECT 233.140000 0.000000 234.830000 0.140000 ;
      RECT 231.240000 0.000000 232.930000 0.140000 ;
      RECT 229.340000 0.000000 231.030000 0.140000 ;
      RECT 227.440000 0.000000 229.130000 0.140000 ;
      RECT 225.540000 0.000000 227.230000 0.140000 ;
      RECT 223.640000 0.000000 225.330000 0.140000 ;
      RECT 221.740000 0.000000 223.430000 0.140000 ;
      RECT 219.840000 0.000000 221.530000 0.140000 ;
      RECT 217.940000 0.000000 219.630000 0.140000 ;
      RECT 216.040000 0.000000 217.730000 0.140000 ;
      RECT 214.140000 0.000000 215.830000 0.140000 ;
      RECT 212.240000 0.000000 213.930000 0.140000 ;
      RECT 210.340000 0.000000 212.030000 0.140000 ;
      RECT 208.440000 0.000000 210.130000 0.140000 ;
      RECT 206.540000 0.000000 208.230000 0.140000 ;
      RECT 204.640000 0.000000 206.330000 0.140000 ;
      RECT 202.740000 0.000000 204.430000 0.140000 ;
      RECT 200.840000 0.000000 202.530000 0.140000 ;
      RECT 198.940000 0.000000 200.630000 0.140000 ;
      RECT 197.040000 0.000000 198.730000 0.140000 ;
      RECT 195.140000 0.000000 196.830000 0.140000 ;
      RECT 193.240000 0.000000 194.930000 0.140000 ;
      RECT 191.340000 0.000000 193.030000 0.140000 ;
      RECT 189.440000 0.000000 191.130000 0.140000 ;
      RECT 187.540000 0.000000 189.230000 0.140000 ;
      RECT 185.640000 0.000000 187.330000 0.140000 ;
      RECT 183.740000 0.000000 185.430000 0.140000 ;
      RECT 181.840000 0.000000 183.530000 0.140000 ;
      RECT 179.940000 0.000000 181.630000 0.140000 ;
      RECT 178.040000 0.000000 179.730000 0.140000 ;
      RECT 176.140000 0.000000 177.830000 0.140000 ;
      RECT 174.240000 0.000000 175.930000 0.140000 ;
      RECT 172.340000 0.000000 174.030000 0.140000 ;
      RECT 170.440000 0.000000 172.130000 0.140000 ;
      RECT 168.540000 0.000000 170.230000 0.140000 ;
      RECT 166.640000 0.000000 168.330000 0.140000 ;
      RECT 164.740000 0.000000 166.430000 0.140000 ;
      RECT 162.840000 0.000000 164.530000 0.140000 ;
      RECT 160.940000 0.000000 162.630000 0.140000 ;
      RECT 159.040000 0.000000 160.730000 0.140000 ;
      RECT 157.140000 0.000000 158.830000 0.140000 ;
      RECT 155.240000 0.000000 156.930000 0.140000 ;
      RECT 153.340000 0.000000 155.030000 0.140000 ;
      RECT 151.440000 0.000000 153.130000 0.140000 ;
      RECT 149.540000 0.000000 151.230000 0.140000 ;
      RECT 147.640000 0.000000 149.330000 0.140000 ;
      RECT 145.740000 0.000000 147.430000 0.140000 ;
      RECT 143.840000 0.000000 145.530000 0.140000 ;
      RECT 141.940000 0.000000 143.630000 0.140000 ;
      RECT 140.040000 0.000000 141.730000 0.140000 ;
      RECT 138.140000 0.000000 139.830000 0.140000 ;
      RECT 136.240000 0.000000 137.930000 0.140000 ;
      RECT 134.340000 0.000000 136.030000 0.140000 ;
      RECT 132.440000 0.000000 134.130000 0.140000 ;
      RECT 130.540000 0.000000 132.230000 0.140000 ;
      RECT 128.640000 0.000000 130.330000 0.140000 ;
      RECT 126.740000 0.000000 128.430000 0.140000 ;
      RECT 124.840000 0.000000 126.530000 0.140000 ;
      RECT 122.940000 0.000000 124.630000 0.140000 ;
      RECT 121.040000 0.000000 122.730000 0.140000 ;
      RECT 119.140000 0.000000 120.830000 0.140000 ;
      RECT 117.240000 0.000000 118.930000 0.140000 ;
      RECT 115.340000 0.000000 117.030000 0.140000 ;
      RECT 113.440000 0.000000 115.130000 0.140000 ;
      RECT 111.540000 0.000000 113.230000 0.140000 ;
      RECT 109.640000 0.000000 111.330000 0.140000 ;
      RECT 107.740000 0.000000 109.430000 0.140000 ;
      RECT 105.840000 0.000000 107.530000 0.140000 ;
      RECT 103.940000 0.000000 105.630000 0.140000 ;
      RECT 102.040000 0.000000 103.730000 0.140000 ;
      RECT 100.140000 0.000000 101.830000 0.140000 ;
      RECT 98.240000 0.000000 99.930000 0.140000 ;
      RECT 96.340000 0.000000 98.030000 0.140000 ;
      RECT 94.440000 0.000000 96.130000 0.140000 ;
      RECT 92.540000 0.000000 94.230000 0.140000 ;
      RECT 90.640000 0.000000 92.330000 0.140000 ;
      RECT 88.740000 0.000000 90.430000 0.140000 ;
      RECT 86.840000 0.000000 88.530000 0.140000 ;
      RECT 84.940000 0.000000 86.630000 0.140000 ;
      RECT 83.040000 0.000000 84.730000 0.140000 ;
      RECT 81.140000 0.000000 82.830000 0.140000 ;
      RECT 79.240000 0.000000 80.930000 0.140000 ;
      RECT 77.340000 0.000000 79.030000 0.140000 ;
      RECT 75.440000 0.000000 77.130000 0.140000 ;
      RECT 73.540000 0.000000 75.230000 0.140000 ;
      RECT 71.640000 0.000000 73.330000 0.140000 ;
      RECT 69.740000 0.000000 71.430000 0.140000 ;
      RECT 67.840000 0.000000 69.530000 0.140000 ;
      RECT 65.940000 0.000000 67.630000 0.140000 ;
      RECT 64.040000 0.000000 65.730000 0.140000 ;
      RECT 62.140000 0.000000 63.830000 0.140000 ;
      RECT 60.240000 0.000000 61.930000 0.140000 ;
      RECT 58.340000 0.000000 60.030000 0.140000 ;
      RECT 56.440000 0.000000 58.130000 0.140000 ;
      RECT 54.540000 0.000000 56.230000 0.140000 ;
      RECT 52.640000 0.000000 54.330000 0.140000 ;
      RECT 50.740000 0.000000 52.430000 0.140000 ;
      RECT 48.840000 0.000000 50.530000 0.140000 ;
      RECT 46.940000 0.000000 48.630000 0.140000 ;
      RECT 45.040000 0.000000 46.730000 0.140000 ;
      RECT 43.140000 0.000000 44.830000 0.140000 ;
      RECT 41.240000 0.000000 42.930000 0.140000 ;
      RECT 39.340000 0.000000 41.030000 0.140000 ;
      RECT 37.440000 0.000000 39.130000 0.140000 ;
      RECT 35.540000 0.000000 37.230000 0.140000 ;
      RECT 33.640000 0.000000 35.330000 0.140000 ;
      RECT 31.740000 0.000000 33.430000 0.140000 ;
      RECT 29.840000 0.000000 31.530000 0.140000 ;
      RECT 27.940000 0.000000 29.630000 0.140000 ;
      RECT 26.040000 0.000000 27.730000 0.140000 ;
      RECT 24.140000 0.000000 25.830000 0.140000 ;
      RECT 22.240000 0.000000 23.930000 0.140000 ;
      RECT 20.340000 0.000000 22.030000 0.140000 ;
      RECT 18.440000 0.000000 20.130000 0.140000 ;
      RECT 16.540000 0.000000 18.230000 0.140000 ;
      RECT 14.640000 0.000000 16.330000 0.140000 ;
      RECT 12.740000 0.000000 14.430000 0.140000 ;
      RECT 10.840000 0.000000 12.530000 0.140000 ;
      RECT 8.940000 0.000000 10.630000 0.140000 ;
      RECT 7.040000 0.000000 8.730000 0.140000 ;
      RECT 5.140000 0.000000 6.830000 0.140000 ;
      RECT 3.240000 0.000000 4.930000 0.140000 ;
      RECT 0.000000 0.000000 3.030000 0.140000 ;
    LAYER metal3 ;
      RECT 0.000000 0.000000 251.180000 248.920000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 251.180000 248.920000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 251.180000 248.920000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 251.180000 248.920000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 251.180000 248.920000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 251.180000 248.920000 ;
    LAYER metal9 ;
      RECT 0.000000 0.000000 251.180000 248.920000 ;
    LAYER metal10 ;
      RECT 0.000000 0.000000 251.180000 248.920000 ;
  END
END aes128key

END LIBRARY
